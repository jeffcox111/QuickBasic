�A|  HL 3           ����������������������������������������        ���������Ѐ        ����������        �����������        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������|       �|       ~|������������������       ���      }���������������������      ���      {����������������������      ���      {����������������������      ���      w����������������������      ���      w���������������������      ����     w���������������������      ����     w��?�������������������      ����     w��?����������������� ��  0������  0{��>r�������������������  0������  0{��>rs����������������������������y�>>rrs�������������������0��������0z|~>rrrs��������������~����0��������0y��>rrrs�������������������0��������0|��~r�������������������<��������<|�������������������      ����     ~?�������������������?�      ���      ��������������������      ���      ���������������������      ��      �������������������        �?�      �������������������        ��      ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ��������������������        �        ����������        �        �        ����������        �        �                  ������������������������������                                                                            