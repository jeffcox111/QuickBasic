�Q�        ���������   � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    � � �    ���������     ���������   � Ȁ � �   �� ��   �� ��   �Ȁ ��   ��� ��   ��� ��   �� �   �� �   �<� �<   �|� �|   �x� �x   ��� ��   ��� ��   ��� ��   ��� ��   ��� ��   ��� ��   � � �    � � �    ���������