��  HL 3           ����������������������������������������        �        0�        ����������        �        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        �������������������        p��      �������������������        p�?�      �������������������        p��       �������������������      p���      ~��������������������      p���      |������������������?�      p����     |?�������������������      p����     x?�?������������������      p����     x�?�������������������      p����     x�?�������������������      p����     x�?������������������� >`  p����>`  x�?������������������� c`  p����c`  x�?������������������� c~>c?p����c~>c?x?�?������������������ cccp����ccc|?������������������� ccccp����cccc|������������������?� ccccp����cccc~�������������������� c~>?p��� c~>? �������������������      p���      �������������������        p��      �������������������        p�?�      �������������������        p��      ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ��������������������        p�        ����������        �����������        ����������        �����������                  ������������������������������                                                                            